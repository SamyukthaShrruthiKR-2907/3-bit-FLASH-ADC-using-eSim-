module samyuktha_flashadc(c,a,b);
input a,b;
output c;
xor (c,a,b);
endmodule